   -- 20ns CLOCK
   --clk <= not clk after 10 ns;