------------------------------


------------------------------