library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package gpu_pkg is
    type array_t is array (0 to 4) of STD_LOGIC_VECTOR(15 downto 0);
end package gpu_pkg;
